library verilog;
use verilog.vl_types.all;
entity divi_freq_vlg_vec_tst is
end divi_freq_vlg_vec_tst;
