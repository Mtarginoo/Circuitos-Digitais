library verilog;
use verilog.vl_types.all;
entity divi_freq_vlg_check_tst is
    port(
        clock_out       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end divi_freq_vlg_check_tst;
