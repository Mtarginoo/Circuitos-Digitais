library verilog;
use verilog.vl_types.all;
entity Dec7Seg_vlg_vec_tst is
end Dec7Seg_vlg_vec_tst;
